`include "../test/core0_base.sv"

module core0_test1;

  initial begin

  end
endmodule
