`define F_DATA_STACK_OVERFLOW 3'h0
`define F_SIGNED_DIVIDE_BY_ZERO 3'h1
`define F_UNSIGNED_DIVIDE_BY_ZERO 3'h2
`define F_SEGFAULT 3'h3
`define F_NONE 3'h7
