`define I_RREADZ 8'b000000ZZ
`define I_RREAD0 8'h00
`define I_RREAD1 8'h01
`define I_RREAD2 8'h02
`define I_RREAD3 8'h03
`define I_ADDZ 8'b000001ZZ
`define I_ADD0 8'h04
`define I_ADD1 8'h05
`define I_ADD2 8'h06
`define I_ADD3 8'h07
`define I_INC 8'h08
`define I_DEC 8'h09
`define I_CARRY 8'h0A
`define I_BORROW 8'h0B
`define I_INV 8'h0C
`define I_BREAK 8'h0D
`define I_READS 8'h0E
`define I_RET 8'h0F
`define I_CONTINUE 8'h10
`define I_IEN 8'h11
`define I_RECV 8'h12
`define I_LD0I 8'h13
`define I_KILL 8'h14
`define I_WAIT 8'h15
`define I_GETBP 8'h16
`define I_GETBA 8'h17
`define I_CALLI 8'h18
`define I_JMPI 8'h19
`define I_JC 8'h1A
`define I_JNC 8'h1B
`define I_JO 8'h1C
`define I_JNO 8'h1D
`define I_JI 8'h1E
`define I_JNI 8'h1F
`define I_CVZ 8'b0010ZZZZ
`define I_READZ 8'b001100ZZ
`define I_READ0 8'h30
`define I_READ1 8'h31
`define I_READ2 8'h32
`define I_READ3 8'h33
`define I_GETZ 8'b001101ZZ
`define I_GET0 8'h34
`define I_GET1 8'h35
`define I_GET2 8'h36
`define I_GET3 8'h37
`define I_IZ 8'b001110ZZ
`define I_I0 8'h38
`define I_I1 8'h39
`define I_I2 8'h3A
`define I_I3 8'h3B
`define I_P0 8'h3C
`define I_READI 8'h3D
`define I_GETP 8'h3E
`define I_GETA 8'h3F
`define I_WRITEZ 8'b010000ZZ
`define I_WRITE0 8'h40
`define I_WRITE1 8'h41
`define I_WRITE2 8'h42
`define I_WRITE3 8'h43
`define I_SETFZ 8'b010001ZZ
`define I_SETF0 8'h44
`define I_SETF1 8'h45
`define I_SETF2 8'h46
`define I_SETF3 8'h47
`define I_SETBZ 8'b010010ZZ
`define I_SETB0 8'h48
`define I_SETB1 8'h49
`define I_SETB2 8'h4A
`define I_SETB3 8'h4B
`define I_ADD 8'h4C
`define I_SUB 8'h4D
`define I_LSL 8'h4E
`define I_LSR 8'h4F
`define I_CSL 8'h50
`define I_CSR 8'h51
`define I_ASR 8'h52
`define I_AND 8'h53
`define I_OR 8'h54
`define I_XOR 8'h55
`define I_READA 8'h56
`define I_CALL 8'h57
`define I_JMP 8'h58
`define I_ISET 8'h59
`define I_SEB 8'h5C
`define I_SLB 8'h5B
`define I_USB 8'h5C
`define I_SEND 8'h5D
`define I_LOOPI 8'h5F
`define I_RAWRITEZ 8'b011000ZZ
`define I_REWRITEZ 8'b011001ZZ
`define I_RAWRITE0 8'h60
`define I_RAWRITE1 8'h61
`define I_RAWRITE2 8'h62
`define I_REWRITE3 8'h63
`define I_REWRITE0 8'h64
`define I_REWRITE1 8'h65
`define I_REWRITE2 8'h66
`define I_REWRITE3 8'h67
`define I_WRITE 8'h68
`define I_WRITEP 8'h69
`define I_WRITEPI 8'h6A
`define I_JEQ 8'h6B
`define I_JNE 8'h6C
`define I_LES 8'h6D
`define I_LEQ 8'h6E
`define I_LESU 8'h6F
`define I_LEQU 8'h70
`define I_IN 8'h71
`define I_OUT 8'h72
`define I_INCEPT 8'h73
`define I_SET 8'h74
`define I_SEL 8'h75
`define I_SETA 8'h76
`define I_LOOP 8'h77
`define I_SEF 8'h78
`define I_MUL 8'h79
`define I_MULU 8'h7A
`define I_DIV 8'h7B
`define I_DIVU 8'h7C
`define I_ROTZ 8'b10ZZZZZZ
`define I_COPYZ 8'b11ZZZZZZ
