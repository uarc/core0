`define OP_LSL 3'h0
`define OP_LSR 3'h1
`define OP_CSL 3'h2
`define OP_CSR 3'h3
`define OP_ASR 3'h4
`define OP_AND 3'h5
`define OP_OR 3'h6
`define OP_ADD 3'h7
