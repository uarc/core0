`define F_DATA_STACK_OVERFLOW 2'h0
`define F_SIGNED_DIVIDE_BY_ZERO 2'h1
`define F_UNSIGNED_DIVIDE_BY_ZERO 2'h2
`define F_SEGFAULT 2'h3
