module core0();

endmodule
